
module reset_ff #(parameter WIDTH = 8) (
    input       clk, rst,
    input       stall,                
    input  [WIDTH-1:0] d,
    output reg [WIDTH-1:0] q
);

always @(posedge clk or posedge rst) begin
    if (rst)
        q <= 0;
    else if (!stall)                  
        q <= d;
 
end

endmodule
